`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05/21/2021 11:52:06 AM
// Design Name: 
// Module Name: noisy
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module noisy(
    input clk,
    input rst_n,

    input signed [13:0] sigin,
    output reg signed [13:0] sigout
    );

    
endmodule
